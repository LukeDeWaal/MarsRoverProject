library IEEE;
use IEEE.std_logic_1164.all;


entity mux_8bit_4input_4sel is
	port (	input_0	: in	std_logic_vector (7 downto 0);
		input_1	: in	std_logic_vector (7 downto 0);
		input_2	: in	std_logic_vector (7 downto 0);
		input_3	: in	std_logic_vector (7 downto 0);
		sel	: in	std_logic_vector (3 downto 0);
		output	: out	std_logic_vector (7 downto 0)
	);
end entity mux_8bit_4input_4sel;

architecture behavioural of mux_8bit_4input_4sel is
begin

	process (input_0, input_1, input_2, input_3, sel)
	begin
		case sel is
			when "1000"	=> output <= input_0;
			when "0100"	=> output <= input_1;
			when "0010"	=> output <= input_2;
			when "0001"	=> output <= input_3;
			when others	=> output <= "00000000";
		end case;
	end process;

end architecture behavioural;
